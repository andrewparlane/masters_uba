library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.fp_type_pkg.all;

entity fp_unpack is
    generic (TBITS:     natural;
             EBITS:     natural);
end entity fp_unpack;

architecture synth of fp_unpack is

begin
end architecture synth;
